--=============================================================================
--Library Declarations:
--=============================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use ieee.math_real.all;
library UNISIM;
use UNISIM.VComponents.all;

--=============================================================================
--Entity Declaration:
--=============================================================================
entity FinalProject_Display is
  Port ( 
      --timing:
    clk_port 	        : in std_logic;
    take_sample_port : in std_logic;
    
    --outputs
    led1 : out std_logic;
    light_output : in std_logic_vector (15 downto 0);
    light_3_bits: out std_logic_vector (2 downto 0);
    led2 : out std_logic;
    led3 : out std_logic;
    led4 : out std_logic;
    led5 : out std_logic);

    
end FinalProject_Display;

--=============================================================================
--Architecture Type:
--=============================================================================
architecture Behavioral of FinalProject_Display is
type state is (NONE,L1,L2,L3,L4,L5);
--=============================================================================
--Signal Declarations: 
    signal current_state, nextState: state := NONE;
    signal light_signal : std_logic_vector (15 downto 0); --4 so that the limit is 15 and each light has 33.3% chance of turning on
    signal mod_value : integer; -- stores a value from 0-4 that corresponds to an LED to turn on 
    signal light_sig_int: integer; -- integer conversion of the number generated by the LFSR
    signal mod_num: integer := 5; --value used to find the mod value 
    constant system_clk_period : time := 10ns;

--=============================================================================



--=============================================================================
--Processes: 
--============================================
--=================================
begin

--state update process
  StateUpdate: process(clk_port,take_sample_port)
  begin
      if rising_edge(clk_port) then 
        if take_sample_port ='1' then
          current_state <= nextState;
          end if;
      end if;

  end process StateUpdate;
  
  NextStateLogic: process(current_state,light_output, light_sig_int,mod_value, mod_num,take_sample_port)
  begin
	nextState <= current_state;
    light_sig_int <= to_integer(signed(light_output));
    mod_value <= light_sig_int mod mod_num;
    
    case current_state is 
   
    	when NONE=>
        	if (mod_value = 0 and light_output/="0000000000000000") then
            	nextState <= L1;
            end if;
            if mod_value = 1  then
            	nextState <= L2;
            end if;
            if mod_value = 2  then
            	nextState <= L3;
            end if;
            if mod_value = 3  then
            	nextState <= L4;
            end if;
            if mod_value = 4  then
            	nextState <= L5;
            end if;
            
  
        when L1 =>
        
        	nextState <= NONE;
        when L2 =>
        	nextState <= NONE;
        when L3 =>
        	nextState <= NONE;
        when L4 =>
        	nextState <= NONE;
        when L5 =>
        	nextState <= NONE;
            
            --edge case
        when others =>
        	nextState <= NONE;
      end case;
  end process NextStateLogic;

  OutputLogic: process(current_state,clk_port)
  begin

--everything starts off with not being enabled 

	led1 <= '0';
    led2 <= '0';
    led3 <= '0';
    led4 <= '0';
    led5 <= '0';
    light_3_bits <= "000";
    case current_state is 
    
        when L1 =>
        	led1 <= '1';
        	led2 <= '0';
            led3 <= '0';
            led4 <= '0';
            led5 <= '0';
        	light_3_bits <= "001";

       	
        when L2 =>
        	led2 <= '1';
        	led1 <= '0';
            led3 <= '0';
            led4 <= '0';
            led5 <= '0';
        	light_3_bits <= "010";
        
        when L3 =>
        	led3 <= '1';
        	led2 <= '0';
            led1 <= '0';
            led4 <= '0';
            led5 <= '0';
        	light_3_bits <= "011";
        
        when L4 =>
        	led4 <= '1';
        	led2 <= '0';
            led3 <= '0';
            led1 <= '0';
            led5 <= '0';
        	light_3_bits <= "100";
            
        when L5 =>
        	led5 <= '1';
        	led2 <= '0';
            led3 <= '0';
            led4 <= '0';
            led1 <= '0';
        	light_3_bits <= "101";
            
        when others =>
        	led1 <= '0';
            led2 <= '0';
            led3 <= '0';
            led4 <= '0';
            led5 <= '0';
            light_3_bits <= "000";
        	
     end case;

    
  end process OutputLogic;
				

  
end behavioral;
